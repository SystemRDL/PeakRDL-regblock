begin
    {%- filter indent %}
    {%- block body %}
    {%- endblock %}
    {%- endfilter %}
end
