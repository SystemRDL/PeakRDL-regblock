{%- block body %}
{%- endblock %}
