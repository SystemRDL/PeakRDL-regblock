// TODO: Add a banner
package {{hwif.package_name}};
    {{hwif.get_package_contents()|indent}}
endpackage
