// USER TEMPLATE OVERRIDE
